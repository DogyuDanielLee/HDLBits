module top_module(
  input a,
  input b,
  input c,
  input d,
  output out  
);
  
  assign out = a | (~b & c);
  // assign out = (a | ~b) & (a | c);
  
endmodule
